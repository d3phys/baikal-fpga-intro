`ifndef __CONTROL_VH__
`define __CONTROL_VH__

// ALU operand (LHS) selector
`define CTL_ALUSEL1_WIDTH   2

`define CTL_ALUSEL1_NONE    `CTL_ALUSEL1_WIDTH'bxx
`define CTL_ALUSEL1_SRC1    `CTL_ALUSEL1_WIDTH'b00
`define CTL_ALUSEL1_UIMM    `CTL_ALUSEL1_WIDTH'b01
`define CTL_ALUSEL1_BIMM    `CTL_ALUSEL1_WIDTH'b10
`define CTL_ALUSEL1_JIMM    `CTL_ALUSEL1_WIDTH'b11

// ALU operand (RHS) selector
`define CTL_ALUSEL2_WIDTH   2

`define CTL_ALUSEL2_NONE    `CTL_ALUSEL2_WIDTH'bxx
`define CTL_ALUSEL2_SRC2    `CTL_ALUSEL2_WIDTH'b00
`define CTL_ALUSEL2_IIMM    `CTL_ALUSEL2_WIDTH'b01
`define CTL_ALUSEL2_SIMM    `CTL_ALUSEL2_WIDTH'b10
`define CTL_ALUSEL2_PC      `CTL_ALUSEL2_WIDTH'b11

// Writeback selector
`define CTL_WBSEL_WIDTH     2

`define CTL_WBSEL_NONE      `CTL_WBSEL_WIDTH'bxx
`define CTL_WBSEL_ALU       `CTL_WBSEL_WIDTH'b00
`define CTL_WBSEL_LSU       `CTL_WBSEL_WIDTH'b01
`define CTL_WBSEL_UIMM      `CTL_WBSEL_WIDTH'b10
`define CTL_WBSEL_PCINC     `CTL_WBSEL_WIDTH'b11

`endif // __CONTROL_VH__
